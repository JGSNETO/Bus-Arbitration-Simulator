library verilog;
use verilog.vl_types.all;
entity busSimulator_vlg_vec_tst is
end busSimulator_vlg_vec_tst;
